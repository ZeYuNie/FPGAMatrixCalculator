`timescale 1ns / 1ps

import matrix_op_selector_pkg::*;
import matrix_op_defs_pkg::*;

module matrix_op_executor_tb;

    // Parameters
    parameter BLOCK_SIZE = 1152;
    parameter ADDR_WIDTH = 14;
    parameter DATA_WIDTH = 32;

    // Signals
    logic clk;
    logic rst_n;
    logic start;
    calc_type_t op_type;
    logic [2:0] matrix_a_id;
    logic [2:0] matrix_b_id;
    logic [31:0] scalar_in;
    logic busy;
    logic done;

    // BRAM Interface (DUT <-> Storage Manager)
    logic [ADDR_WIDTH-1:0] bram_read_addr;
    logic [DATA_WIDTH-1:0] bram_read_data;

    // Storage Manager Interface (DUT Output)
    logic        dut_write_request;
    logic        dut_write_ready;
    logic [2:0]  dut_write_matrix_id;
    logic [7:0]  dut_write_rows;
    logic [7:0]  dut_write_cols;
    logic [7:0]  dut_write_name [0:7];
    logic [DATA_WIDTH-1:0] dut_write_data;
    logic        dut_write_data_valid;
    logic        dut_write_done;
    logic        dut_writer_ready;

    // TB Write Interface (for initialization)
    logic        tb_write_request;
    logic [2:0]  tb_write_matrix_id;
    logic [7:0]  tb_write_rows;
    logic [7:0]  tb_write_cols;
    logic [7:0]  tb_write_name [0:7];
    logic [DATA_WIDTH-1:0] tb_write_data;
    logic        tb_write_data_valid;
    
    // Muxed Signals to Storage Manager
    logic        mux_write_request;
    logic [2:0]  mux_write_matrix_id;
    logic [7:0]  mux_write_rows;
    logic [7:0]  mux_write_cols;
    logic [7:0]  mux_write_name [0:7];
    logic [DATA_WIDTH-1:0] mux_write_data;
    logic        mux_write_data_valid;
    
    // Storage Manager Outputs (Common)
    logic        sm_write_ready;
    logic        sm_write_done;
    logic        sm_writer_ready;

    // Control for Mux
    logic        tb_driving_storage;

    // Clear Interface (Unused)
    logic        clear_request;
    logic        clear_done;
    logic [2:0]  clear_matrix_id;

    assign clear_request = 1'b0;
    assign clear_matrix_id = 3'd0;

    // -------------------------------------------------------------------------
    // Signal Multiplexing
    // -------------------------------------------------------------------------
    always_comb begin
        if (tb_driving_storage) begin
            mux_write_request    = tb_write_request;
            mux_write_matrix_id  = tb_write_matrix_id;
            mux_write_rows       = tb_write_rows;
            mux_write_cols       = tb_write_cols;
            mux_write_name       = tb_write_name;
            mux_write_data       = tb_write_data;
            mux_write_data_valid = tb_write_data_valid;
            
            // Feedback to DUT (hold it off if it tries to write while TB is driving, though shouldn't happen)
            dut_write_ready      = 1'b0;
            dut_writer_ready     = 1'b0;
            dut_write_done       = 1'b0;
        end else begin
            mux_write_request    = dut_write_request;
            mux_write_matrix_id  = dut_write_matrix_id;
            mux_write_rows       = dut_write_rows;
            mux_write_cols       = dut_write_cols;
            mux_write_name       = dut_write_name;
            mux_write_data       = dut_write_data;
            mux_write_data_valid = dut_write_data_valid;
            
            // Feedback from SM to DUT
            dut_write_ready      = sm_write_ready;
            dut_writer_ready     = sm_writer_ready;
            dut_write_done       = sm_write_done;
        end
    end

    // -------------------------------------------------------------------------
    // DUT Instantiation
    // -------------------------------------------------------------------------
    matrix_op_executor #(
        .BLOCK_SIZE(BLOCK_SIZE),
        .ADDR_WIDTH(ADDR_WIDTH),
        .DATA_WIDTH(DATA_WIDTH)
    ) dut (
        .clk                (clk),
        .rst_n              (rst_n),
        .start              (start),
        .op_type            (op_type),
        .matrix_a           (matrix_a_id),
        .matrix_b           (matrix_b_id),
        .scalar_in          (scalar_in),
        .busy               (busy),
        .done               (done),
        .bram_read_addr     (bram_read_addr),
        .bram_data_out      (bram_read_data),
        .write_request      (dut_write_request),
        .write_ready        (dut_write_ready),
        .write_matrix_id    (dut_write_matrix_id),
        .write_rows         (dut_write_rows),
        .write_cols         (dut_write_cols),
        .write_name         (dut_write_name),
        .write_data         (dut_write_data),
        .write_data_valid   (dut_write_data_valid),
        .write_done         (dut_write_done),
        .writer_ready       (dut_writer_ready)
    );

    // -------------------------------------------------------------------------
    // Matrix Storage Manager Instantiation (Real BRAM)
    // -------------------------------------------------------------------------
    matrix_storage_manager #(
        .BLOCK_SIZE(BLOCK_SIZE),
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH),
        .DEPTH(8192 + 1024)
    ) u_storage_manager (
        .clk                (clk),
        .rst_n              (rst_n),
        
        .write_request      (mux_write_request),
        .write_ready        (sm_write_ready),
        .matrix_id          (mux_write_matrix_id),
        .actual_rows        (mux_write_rows),
        .actual_cols        (mux_write_cols),
        .matrix_name        (mux_write_name),
        .data_in            (mux_write_data),
        .data_valid         (mux_write_data_valid),
        .write_done         (sm_write_done),
        .writer_ready       (sm_writer_ready),
        
        .clear_request      (clear_request),
        .clear_done         (clear_done),
        .clear_matrix_id    (clear_matrix_id),
        
        .read_addr          (bram_read_addr),
        .data_out           (bram_read_data)
    );

    // -------------------------------------------------------------------------
    // Clock Generation
    // -------------------------------------------------------------------------
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // -------------------------------------------------------------------------
    // Helper Task: Write Matrix to BRAM
    // -------------------------------------------------------------------------
    task write_matrix_to_bram(
        input logic [2:0] id,
        input logic [7:0] rows,
        input logic [7:0] cols,
        input int         start_val,
        input int         step_val
    );
        int i;
        begin
            tb_driving_storage = 1;
            @(posedge clk);
            
            // Initiate Write Request
            tb_write_request <= 1'b1;
            tb_write_matrix_id <= id;
            tb_write_rows <= rows;
            tb_write_cols <= cols;
            for(int k=0; k<8; k++) tb_write_name[k] <= 8'h41; // 'A'

            // Wait for write_ready
            wait(sm_write_ready);
            @(posedge clk);
            
            // Wait for writer_ready
            wait(sm_writer_ready);
            @(posedge clk);
            
            // Send Data
            for (i = 0; i < rows * cols; i++) begin
                tb_write_data_valid <= 1'b1;
                tb_write_data <= start_val + i * step_val;
                @(posedge clk);
                // Wait if writer becomes not ready
                while (!sm_writer_ready) @(posedge clk);
            end
            
            tb_write_data_valid <= 1'b0;
            tb_write_request <= 1'b0;
            
            // Wait for write_done
            wait(sm_write_done);
            @(posedge clk);
            
            tb_driving_storage = 0;
            @(posedge clk);
        end
    endtask

    // -------------------------------------------------------------------------
    // Debug Monitor
    // -------------------------------------------------------------------------
    initial begin
        forever begin
            @(posedge clk);
            if (start) $display("[%0t] START asserted. Op: %0d", $time, op_type);
            if (done) $display("[%0t] DONE asserted", $time);
            
            // Monitor State Changes (Accessing internal signal)
            // Note: This requires the simulator to support hierarchical access
            // $display("[%0t] State: %0d", $time, dut.state);
        end
    end

    // -------------------------------------------------------------------------
    // Test Sequence
    // -------------------------------------------------------------------------
    initial begin
        // Initialize
        rst_n = 0;
        start = 0;
        op_type = CALC_ADD;
        matrix_a_id = 0;
        matrix_b_id = 0;
        scalar_in = 0;
        
        tb_driving_storage = 0;
        tb_write_request = 0;
        tb_write_data_valid = 0;

        // Reset
        #20 rst_n = 1;
        #20;

        // -------------------------------------------------------
        // Initialize Input Matrices
        // -------------------------------------------------------
        $display("[%0t] Initializing Matrices in BRAM...", $time);
        
        // Matrix 1 (A): 2x2, [[1, 2], [3, 4]]
        write_matrix_to_bram(1, 2, 2, 1, 1);
        
        // Matrix 2 (B): 2x2, [[5, 6], [7, 8]]
        write_matrix_to_bram(2, 2, 2, 5, 1);
        
        $display("[%0t] Initialization Done.", $time);
        #20;

        // -------------------------------------------------------
        // Test 1: Scalar Multiplication
        // -------------------------------------------------------
        $display("[%0t] Test 1: Scalar Multiplication Start", $time);
        op_type = CALC_SCALAR_MUL;
        matrix_a_id = 1; // Use Matrix 1
        scalar_in = 10;  // Scalar = 10
        start = 1;
        #10 start = 0;

        // Wait for completion with timeout
        fork
            begin
                wait(done == 1);
                $display("[%0t] Test 1 Done", $time);
            end
            begin
                #100000; // 100us timeout
                $display("[%0t] Test 1 Timeout! DUT State: %0d", $time, dut.state);
                $finish;
            end
        join_any
        disable fork;
        
        #20;
        
        // Note: Result is in Matrix 0 (ANS).
        // We could verify it by reading BRAM, but for now we trust the done signal
        // and the fact that the simulation didn't hang.
        // Expected: [[10, 20], [30, 40]]

        // -------------------------------------------------------
        // Test 2: Matrix Addition
        // -------------------------------------------------------
        $display("[%0t] Test 2: Matrix Addition Start", $time);
        op_type = CALC_ADD;
        matrix_a_id = 1; // Matrix 1
        matrix_b_id = 2; // Matrix 2
        start = 1;
        #10 start = 0;
        
        fork
            begin
                wait(done == 1);
                $display("[%0t] Test 2 Done", $time);
            end
            begin
                #100000; // 100us timeout
                $display("[%0t] Test 2 Timeout! DUT State: %0d", $time, dut.state);
                $finish;
            end
        join_any
        disable fork;

        #20;
        // Expected: [[6, 8], [10, 12]]

        // -------------------------------------------------------
        // Test 3: Matrix Transpose
        // -------------------------------------------------------
        $display("[%0t] Test 3: Matrix Transpose Start", $time);
        op_type = CALC_TRANSPOSE;
        matrix_a_id = 1; // Matrix 1
        start = 1;
        #10 start = 0;
        
        fork
            begin
                wait(done == 1);
                $display("[%0t] Test 3 Done", $time);
            end
            begin
                #100000; // 100us timeout
                $display("[%0t] Test 3 Timeout! DUT State: %0d", $time, dut.state);
                $finish;
            end
        join_any
        disable fork;

        #20;
        // Expected: [[1, 3], [2, 4]]

        // -------------------------------------------------------
        // Test 4: Convolution
        // -------------------------------------------------------
        $display("[%0t] Test 4: Convolution Start", $time);
        
        // Initialize Matrix 3 (Kernel): 3x3, 1 to 9
        write_matrix_to_bram(3, 3, 3, 1, 1);
        
        op_type = CALC_CONV;
        matrix_a_id = 3; // Matrix 3 (Kernel)
        start = 1;
        #10 start = 0;
        
        fork
            begin
                wait(done == 1);
                $display("[%0t] Test 4 Done", $time);
            end
            begin
                #200000; // 200us timeout (convolution takes longer)
                $display("[%0t] Test 4 Timeout! DUT State: %0d", $time, dut.state);
                $finish;
            end
        join_any
        disable fork;

        #20;

        $display("[%0t] All Tests Passed", $time);
        $finish;
    end

endmodule
