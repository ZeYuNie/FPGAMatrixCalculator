`timescale 1ps / 1ps

module settings_ram (
    input  logic         clk,
    input  logic         rst_n,

    input  logic         valid_set_max_row,
    input  logic         valid_set_max_col,
    input  logic         valid_data_min,
    input  logic         valid_data_max,

    input  

)